  parameter zero = 'b00111111;
  parameter um = 'b00000110;
  parameter dois = 'b01011011;
  parameter tres = 'b01001111;
  parameter quatro = 'b01100110;
  parameter cinco = 'b01101101;
  parameter seis = 'b01111101;
  parameter sete = 'b00000111;
  parameter oito = 'b01111111;
  parameter nove = 'b01101111;
  parameter dez = 'b01110111;
  parameter onze = 'b01111111;
  parameter doze = 'b00111001;
  parameter treze = 'b00111111;
  parameter quatorze = 'b01111001;
  parameter quinze = 'b01110001;

  parameter Lzero = 'b0000;
  parameter Lum = 'b0001;
  parameter Ldois = 'b0010;
  parameter Ltres = 'b0011;
  parameter Lquatro = 'b0100;
  parameter Lcinco = 'b0101;
  parameter Lseis = 'b0110;
  parameter Lsete = 'b0111;
  parameter Loito = 'b1000;
  parameter Lnove = 'b1001;
  parameter Ldez = 'b1010;
  parameter Lonze = 'b1011;
  parameter Ldoze = 'b1100;
  parameter Ltreze = 'b1101;
  parameter Lquatorze = 'b1110;
  parameter Lquinze = 'b1111;